module multiplexer_2_1(
	input a,
	input b,
	input select,
	output y
);
	assign y = (select)?b:a;
endmodule
